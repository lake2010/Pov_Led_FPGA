library verilog;
use verilog.vl_types.all;
entity Qsys_system_mm_interconnect_0 is
    port(
        clk_clk_clk     : in     vl_logic;
        nios2_qsys_reset_n_reset_bridge_in_reset_reset: in     vl_logic;
        nios2_qsys_data_master_address: in     vl_logic_vector(15 downto 0);
        nios2_qsys_data_master_waitrequest: out    vl_logic;
        nios2_qsys_data_master_byteenable: in     vl_logic_vector(3 downto 0);
        nios2_qsys_data_master_read: in     vl_logic;
        nios2_qsys_data_master_readdata: out    vl_logic_vector(31 downto 0);
        nios2_qsys_data_master_readdatavalid: out    vl_logic;
        nios2_qsys_data_master_write: in     vl_logic;
        nios2_qsys_data_master_writedata: in     vl_logic_vector(31 downto 0);
        nios2_qsys_data_master_debugaccess: in     vl_logic;
        nios2_qsys_instruction_master_address: in     vl_logic_vector(15 downto 0);
        nios2_qsys_instruction_master_waitrequest: out    vl_logic;
        nios2_qsys_instruction_master_read: in     vl_logic;
        nios2_qsys_instruction_master_readdata: out    vl_logic_vector(31 downto 0);
        nios2_qsys_instruction_master_readdatavalid: out    vl_logic;
        epcs_flash_epcs_control_port_address: out    vl_logic_vector(8 downto 0);
        epcs_flash_epcs_control_port_write: out    vl_logic;
        epcs_flash_epcs_control_port_read: out    vl_logic;
        epcs_flash_epcs_control_port_readdata: in     vl_logic_vector(31 downto 0);
        epcs_flash_epcs_control_port_writedata: out    vl_logic_vector(31 downto 0);
        epcs_flash_epcs_control_port_chipselect: out    vl_logic;
        Hal249_s1_address: out    vl_logic_vector(1 downto 0);
        Hal249_s1_write : out    vl_logic;
        Hal249_s1_readdata: in     vl_logic_vector(31 downto 0);
        Hal249_s1_writedata: out    vl_logic_vector(31 downto 0);
        Hal249_s1_chipselect: out    vl_logic;
        jtag_uart_avalon_jtag_slave_address: out    vl_logic_vector(0 downto 0);
        jtag_uart_avalon_jtag_slave_write: out    vl_logic;
        jtag_uart_avalon_jtag_slave_read: out    vl_logic;
        jtag_uart_avalon_jtag_slave_readdata: in     vl_logic_vector(31 downto 0);
        jtag_uart_avalon_jtag_slave_writedata: out    vl_logic_vector(31 downto 0);
        jtag_uart_avalon_jtag_slave_waitrequest: in     vl_logic;
        jtag_uart_avalon_jtag_slave_chipselect: out    vl_logic;
        Led_s1_address  : out    vl_logic_vector(1 downto 0);
        Led_s1_write    : out    vl_logic;
        Led_s1_readdata : in     vl_logic_vector(31 downto 0);
        Led_s1_writedata: out    vl_logic_vector(31 downto 0);
        Led_s1_chipselect: out    vl_logic;
        nios2_qsys_jtag_debug_module_address: out    vl_logic_vector(8 downto 0);
        nios2_qsys_jtag_debug_module_write: out    vl_logic;
        nios2_qsys_jtag_debug_module_read: out    vl_logic;
        nios2_qsys_jtag_debug_module_readdata: in     vl_logic_vector(31 downto 0);
        nios2_qsys_jtag_debug_module_writedata: out    vl_logic_vector(31 downto 0);
        nios2_qsys_jtag_debug_module_byteenable: out    vl_logic_vector(3 downto 0);
        nios2_qsys_jtag_debug_module_waitrequest: in     vl_logic;
        nios2_qsys_jtag_debug_module_debugaccess: out    vl_logic;
        onchip_ram_s1_address: out    vl_logic_vector(11 downto 0);
        onchip_ram_s1_write: out    vl_logic;
        onchip_ram_s1_readdata: in     vl_logic_vector(31 downto 0);
        onchip_ram_s1_writedata: out    vl_logic_vector(31 downto 0);
        onchip_ram_s1_byteenable: out    vl_logic_vector(3 downto 0);
        onchip_ram_s1_chipselect: out    vl_logic;
        onchip_ram_s1_clken: out    vl_logic;
        sysid_qsys_control_slave_address: out    vl_logic_vector(0 downto 0);
        sysid_qsys_control_slave_readdata: in     vl_logic_vector(31 downto 0)
    );
end Qsys_system_mm_interconnect_0;
